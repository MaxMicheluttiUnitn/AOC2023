module main
import partone
import parttwo

fn main() {
	// partone.partone('problem.txt')!
	parttwo.parttwo('problem.txt')!
}
